module DeBounce(clk,reset,button_in,DB_out);
	
input clk,reset,button_in,DB_out;

endmodule


